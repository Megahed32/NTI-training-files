`include "uvm_macros.svh"
`include "interface.sv"

package driver_pkg;

import uvm_pkg::*;
import transaction_pkg::*;

class my_driver extends uvm_driver #(my_sequence_item);

    `uvm_component_utils(my_driver);
        virtual intf vif_driver;
        my_sequence_item seq_item;

    function new(string name = "my_driver" , uvm_component parent = null);
        super.new(name , parent);
    endfunction

    function void build_phase(uvm_phase phase);
        super.build_phase(phase);
        if (!(uvm_config_db #(virtual intf)::get(this , "" , "my_vif" , vif_driver)))
        `uvm_info("Getting VIF in driver", $sformatf("Failed"), UVM_LOW);
        $display("driver build phase");
    endfunction

    function void connect_phase(uvm_phase phase);
        super.connect_phase(phase);
        $display("driver connect phase");
    endfunction

    task run_phase(uvm_phase phase);
        super.run_phase(phase);

        $display("driver run phase");
        forever
        begin
        seq_item_port.get_next_item(seq_item);
        // Drive signals to DUT
        @(negedge vif_driver.clk);
        vif_driver.rst      = seq_item.rst;
        vif_driver.re       = seq_item.re;
        vif_driver.en       = seq_item.en;
        vif_driver.addr     = seq_item.addr;       
        vif_driver.data_in  = seq_item.data_in;
        
        seq_item_port.item_done();
        end 
    endtask
endclass





endpackage